`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/08/06 10:01:06
// Design Name: 
// Module Name: LabMain
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module LabMain(A, clk, rst, AN, Seg);

input [4:0] A;
input clk, rst;
output [7:0] AN;
output [7:0] Seg;

wire [4:0] outbit;

MainBlock U1(.ib(A), .ob(outbit));
Dsp7Seg U2 (.X0(outbit[0]), .X1(outbit[1]), .X2(outbit[2]), .X3(outbit[3]), .X4(outbit[4]), .clk(clk), .rst(rst), .AN(AN), .dsp(Seg));

endmodule
